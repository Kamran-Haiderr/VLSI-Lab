* SPICE netlist written by S-Edit Win32 7.00
* Written on Nov 19, 2001 at 08:40:00

* No Ports in cell: <MacroCalls>
* End of module with no ports: <MacroCalls>

* No Ports in cell: PageID_Tanner
* End of module with no ports: PageID_Tanner

.SUBCKT DFFC ClB Clk Data Q QB Gnd Vdd
MN_4_1 10 4 Gnd Gnd NMOS W='15*l' L='2*l' AS='72*l*l' AD='45*l*l' PS='42*l' PD='21*l' M=1
MN_4_2 14 Q Gnd Gnd NMOS W='22*l' L='2*l' AS='66*l*l' AD='22*l*l' PS='28*l' PD='24*l' M=1
MN_4_3 8 ClB Gnd Gnd NMOS W='15*l' L='2*l' AS='45*l*l' AD='15*l*l' PS='21*l' PD='17*l' M=1
MN_4_4 C CB Gnd Gnd NMOS W='6*l' L='2*l' AS='43.7778*l*l' AD='36*l*l' PS='18.2222*l' PD='24*l' M=1
MN_4_5 CB Clk Gnd Gnd NMOS W='6*l' L='2*l' AS='43.7778*l*l' AD='42*l*l' PS='18.2222*l' PD='26*l' M=1
MN_4_6 Q 12 Gnd Gnd NMOS W='22*l' L='2*l' AS='185*l*l' AD='66*l*l' PS='64*l' PD='28*l' M=1
MN_4_7 12 CB QB Gnd NMOS W='15*l' L='2*l' AS='45*l*l' AD='59.5946*l*l' PS='21*l' PD='23.5135*l' M=1
MN_4_8 QB ClB 14 Gnd NMOS W='22*l' L='2*l' AS='22*l*l' AD='87.4054*l*l' PS='24*l' PD='34.4865*l' M=1
MN_4_9 12 C 13 Gnd NMOS W='15*l' L='2*l' AS='45*l*l' AD='15*l*l' PS='21*l' PD='17*l' M=1
MN_4_10 13 10 Gnd Gnd NMOS W='15*l' L='2*l' AS='15*l*l' AD='123*l*l' PS='17*l' PD='50*l' M=1
MN_4_11 4 C 7 Gnd NMOS W='15*l' L='2*l' AS='45*l*l' AD='45*l*l' PS='21*l' PD='21*l' M=1
MN_4_12 7 10 8 Gnd NMOS W='15*l' L='2*l' AS='15*l*l' AD='45*l*l' PS='17*l' PD='21*l' M=1
MN_4_13 4 CB 5 Gnd NMOS W='15*l' L='2*l' AS='45*l*l' AD='15*l*l' PS='21*l' PD='17*l' M=1
MN_4_14 5 Data Gnd Gnd NMOS W='15*l' L='2*l' AS='15*l*l' AD='109.444*l*l' PS='17*l' PD='45.5556*l' M=1
* Page Size:  5x7
* S-Edit  D Flip-Flop with Clear (TIB)
* Designed by: J. Luo  Jul 17, 1998  12:22:28
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module DFFC / page Page0 
MP_4_1 QB Q Vdd Vdd PMOS W='24*l' L='2*l' AS='114*l*l' AD='72*l*l' PS='60*l' PD='30*l' M=1
MP_4_2 10 4 Vdd Vdd PMOS W='15*l' L='2*l' AS='90*l*l' AD='86.25*l*l' PS='42*l' PD='38.75*l' M=1
MP_4_3 4 CB 9 Vdd PMOS W='11*l' L='2*l' AS='33.55*l*l' AD='47.6667*l*l' PS='18.7*l' PD='18.8571*l' M=1
MP_4_4 9 ClB Vdd Vdd PMOS W='9*l' L='2*l' AS='51.75*l*l' AD='27.45*l*l' PS='23.25*l' PD='15.3*l' M=1
MP_4_5 C CB Vdd Vdd PMOS W='6*l' L='2*l' AS='36*l*l' AD='43.8621*l*l' PS='24*l' PD='16.9655*l' M=1
MP_4_6 CB Clk Vdd Vdd PMOS W='6*l' L='2*l' AS='36*l*l' AD='43.8621*l*l' PS='24*l' PD='16.9655*l' M=1
MP_4_7 Q 12 Vdd Vdd PMOS W='27*l' L='2*l' AS='143*0.000001*l' AD='111*l*l' PS='66*l' PD='66*l' M=1
MP_4_8 QB ClB Vdd Vdd PMOS W='24*l' L='2*l' AS='72*l*l' AD='81.6*l*l' PS='30*l' PD='36*l' M=1
MP_4_9 12 C QB Vdd PMOS W='16*l' L='2*l' AS='54.4*l*l' AD='48*l*l' PS='24*l' PD='22*l' M=1
MP_4_10 11 10 Vdd Vdd PMOS W='16*l' L='2*l' AS='16*l*l' AD='96*l*l' PS='18*l' PD='44*l' M=1
MP_4_11 12 CB 11 Vdd PMOS W='16*l' L='2*l' AS='48*l*l' AD='16*l*l' PS='22*l' PD='18*l' M=1
MP_4_12 6 10 Vdd Vdd PMOS W='14*l' L='2*l' AS='84*l*l' AD='14*l*l' PS='40*l' PD='16*l' M=1
MP_4_13 4 CB 6 Vdd PMOS W='14*l' L='2*l' AS='14*l*l' AD='60.6667*l*l' PS='16*l' PD='24*l' M=1
MP_4_14 3 Data Vdd Vdd PMOS W='17*l' L='2*l' AS='17*l*l' AD='124.276*l*l' PS='19*l' PD='48.069*l' M=1
MP_4_15 4 C 3 Vdd PMOS W='17*l' L='2*l' AS='73.6667*l*l' AD='17*l*l' PS='29.1429*l' PD='19*l' M=1
.ENDS

.SUBCKT NAND2C A B Out1 Out2 Gnd Vdd
MN_4_1 Out2 Out1 Gnd Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='122*l*l' PS='68*l' PD='47*l' M=1
MN_4_2 1 B Gnd Gnd NMOS W='28*l' L='2*l' AS='122*l*l' AD='28*l*l' PS='47*l' PD='30*l' M=1
MN_4_3 Out1 A 1 Gnd NMOS W='28*l' L='2*l' AS='28*l*l' AD='148*l*l' PS='30*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  Traffic Light Controller Example
* Designed by: D.Gunawan, J.Luo  Jul 17, 1998  12:22:28
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module NAND2C / page Page0 
MP_4_1 Out2 Out1 Vdd Vdd PMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
MP_4_2 Out1 B Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
MP_4_3 Out1 A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
.ENDS

.SUBCKT NAND3C A B C Out1 Out2 Gnd Vdd
MN_4_1 Out2 Out1 Gnd Gnd NMOS W='28*l' L='2*l' AS='120*l*l' AD='148*l*l' PS='48*l' PD='68*l' M=1
MN_4_2 2 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='120*l*l' PS='34*l' PD='48*l' M=1
MN_4_3 1 B 2 Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
MN_4_4 Out1 C 1 Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
* Page Size:  5x7
* S-Edit  Traffic Light Controller Example
* Designed by: D.Gunawan, J.Luo  Jul 17, 1998  12:22:29
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module NAND3C / page Page0 
MP_4_1 Out2 Out1 Vdd Vdd PMOS W='28*l' L='2*l' AS='122*l*l' AD='148*l*l' PS='47*l' PD='68*l' M=1
MP_4_2 Out1 C Vdd Vdd PMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
MP_4_3 Out1 B Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
MP_4_4 Out1 A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='122*l*l' PS='34*l' PD='47*l' M=1
.ENDS

.SUBCKT NOR2C A B Out1 Out2 Gnd Vdd
MN_4_1 Out2 Out1 Gnd Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
MN_4_2 Out1 B Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
MN_4_3 Out1 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  Traffic Light Controller Example
* Designed by: D.Gunawan, J.Luo  Jul 17, 1998  12:22:29
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module NOR2C / page Page0 
MP_4_1 Out2 Out1 Vdd Vdd PMOS W='28*l' L='2*l' AS='148*l*l' AD='122*l*l' PS='68*l' PD='47*l' M=1
MP_4_2 Out1 A 1 Vdd PMOS W='28*l' L='2*l' AS='28*l*l' AD='148*l*l' PS='30*l' PD='68*l' M=1
MP_4_3 1 B Vdd Vdd PMOS W='28*l' L='2*l' AS='122*l*l' AD='28*l*l' PS='47*l' PD='30*l' M=1
.ENDS

.SUBCKT NOR2 A B Out Gnd Vdd
MN_4_1 Out B Gnd Gnd NMOS W='28*l' L='2*l' AS='144*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
MN_4_2 Out A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
* Page Size:  5x7
* S-Edit  2-Input NOR Gate (TIB)
* Designed by: J. Luo  Jul 17, 1998  12:22:29
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module NOR2 / page Page0 
MP_4_1 Out B 1 Vdd PMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
MP_4_2 1 A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='144*l*l' PS='34*l' PD='68*l' M=1
.ENDS

.SUBCKT NOR3C A B C Out1 Out2 Gnd Vdd
MN_4_1 Out2 Out1 Gnd Gnd NMOS W='28*l' L='2*l' AS='122*l*l' AD='148*l*l' PS='47*l' PD='68*l' M=1
MN_4_2 Out1 C Gnd Gnd NMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
MN_4_3 Out1 B Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
MN_4_4 Out1 A Gnd Gnd NMOS W='28*l' L='2*l' AS='84*l*l' AD='122*l*l' PS='34*l' PD='47*l' M=1
* Page Size:  5x7
* S-Edit  Traffic Light Controller Example
* Designed by: D.Gunawan, J.Luo  Jul 17, 1998  12:22:29
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module NOR3C / page Page0 
MP_4_1 Out2 Out1 Vdd Vdd PMOS W='28*l' L='2*l' AS='122*l*l' AD='148*l*l' PS='47*l' PD='68*l' M=1
MP_4_2 Out1 C 2 Vdd PMOS W='28*l' L='2*l' AS='148*l*l' AD='84*l*l' PS='68*l' PD='34*l' M=1
MP_4_3 2 B 1 Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='84*l*l' PS='34*l' PD='34*l' M=1
MP_4_4 1 A Vdd Vdd PMOS W='28*l' L='2*l' AS='84*l*l' AD='122*l*l' PS='34*l' PD='47*l' M=1
.ENDS

* No Ports in cell: Page5x7
* End of module with no ports: Page5x7

.SUBCKT core CLOCK DONT_EW DONT_NS GREEN_EW GREEN_NS RED_EW RED_NS RESETB
+ TEST_POINT TOP4 TOP5 TOP6 WALK_EW WALK_NS YELLOW_EW YELLOW_NS Gnd Vdd
XDFFC_1 RESETB CLOCK N1 N22 N1 Gnd Vdd DFFC
XDFFC_2 RESETB N1 N3 N7 N3 Gnd Vdd DFFC
XDFFC_3 RESETB N3 N20 N10 N20 Gnd Vdd DFFC
XDFFC_4 RESETB N20 N6 TOP4 N6 Gnd Vdd DFFC
XDFFC_5 RESETB N6 TEST_POINT TOP5 TEST_POINT Gnd Vdd DFFC
XDFFC_6 RESETB TEST_POINT N2 TOP6 N2 Gnd Vdd DFFC
XDFFC_7 RESETB N2 RED_NS RED_EW RED_NS Gnd Vdd DFFC
XNAND2C_1 N5 RED_EW N8 GREEN_NS Gnd Vdd NAND2C
XNAND2C_2 N5 RED_NS N9 GREEN_EW Gnd Vdd NAND2C
XNAND3C_1 N22 TOP6 TEST_POINT N12 N40 Gnd Vdd NAND3C
XNOR2C_1 TEST_POINT N2 N13 N5 Gnd Vdd NOR2C
XNOR2_2 RED_NS N5 YELLOW_NS Gnd Vdd NOR2
XNOR2_5 RED_NS TOP6 WALK_NS Gnd Vdd NOR2
XNOR2_6 TOP6 RED_EW WALK_EW Gnd Vdd NOR2
XNOR2_7 RED_EW N5 YELLOW_EW Gnd Vdd NOR2
XNOR3C_1 N40 YELLOW_NS RED_NS N11 DONT_NS Gnd Vdd NOR3C
XNOR3C_2 N40 YELLOW_EW RED_EW N4 DONT_EW Gnd Vdd NOR3C
* S-Edit  Traffic Light Controller
* Designed by: Jin Luo, Owen Smith  Apr 26, 1996  12:53:42
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module core / page Page0 
.ENDS

.SUBCKT PadGnd PAD Gnd
C1 Gnd Gnd 0.25pF
* Page Size:  5x7
* S-Edit  Ground Pad
* Designed by: D.Gunawan, J.Luo  Nov 19, 2001  11:59:46
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module PadGnd / page Page0 
.ENDS

* No Ports in cell: Substrate
* End of module with no ports: Substrate

.SUBCKT Pad_Bond SIGNAL Gnd
C1 SIGNAL Gnd 0.25pF
* Page Size:  5x7
* S-Edit  Output Pad
* Designed by: D.Gunawan, J.Luo, K.Schaefer  Nov 14, 2001  09:50:47
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module Pad_Bond / page Page0 
.ENDS

.SUBCKT PadBidirHE_2.0u DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Vdd
MN_4_1 OEB OE Gnd Gnd NMOS W=12u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_2 N2 DataOut Gnd Gnd NMOS W=12u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_3 N1 OE N2 Gnd NMOS W=12u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_4 N2 OEB Gnd Gnd NMOS W=12u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_5 Pad N2 Gnd Gnd NMOS W=14.8u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MN_4_6 DataInB DataInUnBuf Gnd Gnd NMOS W=22u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MN_4_7 DataIn DataInB Gnd Gnd NMOS W=13u L=2u AS=66p AD=66p PS=24u PD=24u M=4
XPad_Bond_1 Pad Gnd Pad_Bond
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Nov 14, 2001  13:56:08
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module PadBidirHE_2.0u / page Page0 
MP_4_1 OEB OE Vdd Vdd PMOS W=13u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_2 N1 DataOut Vdd Vdd PMOS W=13u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_3 N2 OEB N1 Vdd PMOS W=13u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_4 N1 OE Vdd Vdd PMOS W=13u L=2u AS=66p AD=66p PS=24u PD=24u M=1
MP_4_5 Pad N1 Vdd Vdd PMOS W=16u L=2u AS=66p AD=66p PS=24u PD=24u M=10
MP_4_6 DataInB DataInUnBuf Vdd Vdd PMOS W=13u L=2u AS=66p AD=66p PS=24u PD=24u M=2
MP_4_7 DataIn DataInB Vdd Vdd PMOS W=55u L=2u AS=66p AD=66p PS=24u PD=24u M=1
R1 Pad DataInUnBuf 84.2333 TC1=0.0 TC2=0.0
.ENDS

.SUBCKT PadBidirHE DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Vdd
XPadBidirHE_2.0u_1 DataIn DataInB DataInUnBuf DataOut OE Pad Gnd Vdd
+ PadBidirHE_2.0u
* Page Size:  5x7
* S-Edit  Bidirectional Pad
* Designed by: D.Gunawan, J.Luo  Jul 17, 1998  12:22:30
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module PadBidirHE / page Page0 
.ENDS

.SUBCKT PadInC DataIn DataInB DataInUnBuf PAD Gnd Vdd
XPadBidirHE_1 DataIn DataInB DataInUnBuf Gnd Gnd PAD Gnd Vdd PadBidirHE
* Page Size:  5x7
* S-Edit  Input Pad
* Designed by: D.Gunawan, J.Luo  Nov 20, 1998  16:27:59
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module PadInC / page Page0 
.ENDS

.SUBCKT PadOut DataOut PAD Gnd Vdd
XPadBidirHE_N20_1 N3 N2 N1 DataOut Vdd PAD Gnd Vdd PadBidirHE_2.0u
* Page Size:  5x7
* S-Edit  SCMOS Library
* Designed by: D.Gunawan, J.Luo, K.Schaefer  Nov 20, 1998  16:26:23
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module PadOut / page Page0 
.ENDS

.SUBCKT PadVdd PAD Gnd Vdd
C1 Vdd Gnd 0.25pF
* Page Size:  5x7
* S-Edit  Vdd Pad
* Designed by: D.Gunawan, J.Luo  Nov 19, 2001  13:25:13
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module PadVdd / page Page0 
.ENDS

* Main circuit: Lights
.include ext_devc.md
.param l=1u
Xcore_1 N21 N15 N45 N13 N41 N11 N37 N9 N8 N7 N6 N5 N4 N43 N2 N39 Gnd Vdd core
XPadGnd_1 PAD_R3 Gnd PadGnd
XPadInC_1 N21 N20 N19 PAD_L2 Gnd Vdd PadInC
XPadInC_2 N9 N24 N23 PAD_L1 Gnd Vdd PadInC
XPadOut_1 N11 PAD_R1 Gnd Vdd PadOut
XPadOut_2 N2 PAD_B3 Gnd Vdd PadOut
XPadOut_3 N13 PAD_B2 Gnd Vdd PadOut
XPadOut_4 N4 PAD_B1 Gnd Vdd PadOut
XPadOut_5 N15 PAD_L4 Gnd Vdd PadOut
XPadOut_6 N37 PAD_R2 Gnd Vdd PadOut
XPadOut_7 N39 PAD_T3 Gnd Vdd PadOut
XPadOut_8 N41 PAD_T2 Gnd Vdd PadOut
XPadOut_9 N43 PAD_T1 Gnd Vdd PadOut
XPadOut_10 N45 PAD_R4 Gnd Vdd PadOut
XPadVdd_1 PAD_L3 Gnd Vdd PadVdd
* S-Edit  Traffic Light Controller Example
* Designed by: Jin Luo, Owen Smith  Nov 19, 2001  13:24:27
* Schematic generated by S-Edit
* from file C:\Tanner\LEdit84\Samples\SPR\example1\lights_tpr / module Lights / page Page0 
* End of main circuit: Lights
.END
