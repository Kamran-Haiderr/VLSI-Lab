* SPICE netlist written by S-Edit Win32 8.10
* Written on Dec 12, 2003 at 11:55:18

.SUBCKT ALU C0 C1 C2 C3 C4 C5 D0 D1 D2 D3 D4 D5 D6 D7
.ENDS

.SUBCKT BUF CLK IN OUT
.ENDS

.SUBCKT CTRL A0 A1 A2 B0 B1 B2 B3 B4 B5 C0 C1 C2 C4 CLK F0 F1
.ENDS

.SUBCKT IOBUF A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15 B0 B1 B2 B3
+ B4 B5 B6 B7 C0 C1 C2 D0 D1 D2 D3 D4 D5 D6 D7
.ENDS

.SUBCKT IOPAD A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15 CLK D0 D1
+ D2 D3 D4 D5 D6 D7
.ENDS

.SUBCKT PC CLK R0 R1 R2 R3 R4 R5 R6 R7
.ENDS

.SUBCKT REG C0 C1 C2 C4 F0 F1 R0 R1 R2 R3 R4 R5 R6 R7
.ENDS

* Main circuit: CPU
XALU_1 N1 N2 N3 N4 N5 N6 D0 D1 D2 D3 D4 D5 D6 D7 ALU
XBUF_1 CLK N53 N1 BUF
XBUF_2 CLK N54 N2 BUF
XBUF_3 CLK N55 N3 BUF
XBUF_4 CLK N56 N4 BUF
XBUF_5 CLK N57 N5 BUF
XBUF_6 CLK N58 N6 BUF
XCTRL_1 N40 N41 N42 N53 N54 N55 N56 N57 N58 N96 N33 N34 N35 CLK N36 N37 CTRL
XIOBUF_1 N88 N87 N86 N85 N84 N83 N82 N81 N80 N79 N78 N77 N76 N75 N74 N73 N89 N91
+ N90 N93 N92 N95 N94 N38 N40 N41 N42 D0 D1 D2 D3 D4 D5 D6 D7 IOBUF
XIOPAD_1 N88 N87 N86 N85 N84 N83 N82 N81 N80 N79 N78 N77 N76 N75 N74 N73 CLK N89
+ N91 N90 N93 N92 N95 N94 N38 IOPAD
XPC_1 CLK D0 D1 D2 D3 D4 D5 D6 D7 PC
XREG_1 N96 N33 N34 N35 N36 N37 D0 D1 D2 D3 D4 D5 D6 D7 REG
* End of main circuit: CPU
.END
